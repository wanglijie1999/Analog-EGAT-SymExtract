** Generated for: hspiceD
** Generated on: Mar  6 21:53:50 2023
** Design library name: proj_DDA
** Design cell name: test3_4
** Design view name: schematic



** Library name: proj_DDA
** Cell name: test3_4
** View name: schematic
.subckt 09DDAWXN vss vout vdd iss _net0 _net1 _net2 _net3
xm34 vdd vdd vdd vdd pch_5 l=500e-9 w=10e-6 m=4 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm35 vdd vdd vdd vdd pch_5 l=500e-9 w=10e-6 m=4 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm36 net54 net54 net54 net54 pch_5 l=500e-9 w=10e-6 m=4 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm37 net31 net31 net31 net31 pch_5 l=500e-9 w=10e-6 m=4 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm40 vdd vdd vdd vdd pch_5 l=2e-6 w=10e-6 m=1 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm20 net019 net029 net20 vdd pch_5 l=1e-6 w=10e-6 m=1 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm41 vdd vdd vdd vdd pch_5 l=1e-6 w=10e-6 m=1 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm17 net20 net019 vdd vdd pch_5 l=2e-6 w=10e-6 m=1 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm15 net58 net019 vdd vdd pch_5 l=2e-6 w=10e-6 m=10 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm14 net54 net029 net58 vdd pch_5 l=1e-6 w=10e-6 m=10 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm30 net33 _net0 net54 net54 pch_5 l=2e-6 w=10e-6 m=8 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm29 net30 _net2 net54 net54 pch_5 l=2e-6 w=10e-6 m=8 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm28 net40 net029 net41 vdd pch_5 l=1e-6 w=10e-6 m=6 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm21 net59 net019 vdd vdd pch_5 l=2e-6 w=10e-6 m=10 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm32 net30 _net1 net31 net31 pch_5 l=2e-6 w=10e-6 m=8 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm31 net33 _net3 net31 net31 pch_5 l=2e-6 w=10e-6 m=8 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm23 net41 net019 vdd vdd pch_5 l=2e-6 w=10e-6 m=6 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm22 net61 net019 vdd vdd pch_5 l=2e-6 w=10e-6 m=6 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm26 vout net029 net61 vdd pch_5 l=1e-6 w=10e-6 m=6 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm25 net31 net029 net59 vdd pch_5 l=1e-6 w=10e-6 m=10 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm44 vss vss vss vss nch_5 l=600e-9 w=8e-6 m=2 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm38 vss vss vss vss nch_5 l=600e-9 w=10e-6 m=2 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm39 vss vss vss vss nch_5 l=600e-9 w=8e-6 m=2 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm27 net064 net012 vss vss nch_5 l=1e-6 w=8e-6 m=1 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm24 net012 net012 vss vss nch_5 l=1e-6 w=8e-6 m=1 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm42 iss iss net012 vss nch_5 l=1e-6 w=8e-6 m=1 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm43 net029 iss net064 vss nch_5 l=1e-6 w=8e-6 m=1 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm7 net33 net40 vss vss nch_5 l=2e-6 w=8e-6 m=1 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm33 net30 net40 vss vss nch_5 l=2e-6 w=8e-6 m=1 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm5 vout iss net30 vss nch_5 l=2e-6 w=10e-6 m=2 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm4 net40 iss net33 vss nch_5 l=2e-6 w=10e-6 m=2 nf=1 sd=540e-9 ad=4.8e-12 as=4.8e-12 pd=20.96e-6 ps=20.96e-6 nrd=27e-3 nrs=27e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xr1  net019 net019   rppolyhri3d3k lr=7.34e-6 wr=1e-6 mf=1 m=1 mismatchflag=1
xr2  net029 net029   rppolyhri3d3k lr=7.34e-6 wr=1e-6 mf=1 m=1 mismatchflag=1

xr0_1__dmy0  net019 xr0_1__dmy0  rppolyhri3d3k lr=7.34e-6 wr=2e-6 mf=1 m=1 mismatchflag=1
xr0_2__dmy0  xr0_1__dmy0 xr0_2__dmy0  rppolyhri3d3k lr=7.34e-6 wr=2e-6 mf=1 m=1 mismatchflag=1
xr0_3__dmy0  xr0_2__dmy0 xr0_3__dmy0  rppolyhri3d3k lr=7.34e-6 wr=2e-6 mf=1 m=1 mismatchflag=1
xr0_4__dmy0  xr0_3__dmy0 xr0_4__dmy0  rppolyhri3d3k lr=7.34e-6 wr=2e-6 mf=1 m=1 mismatchflag=1
xr0_5__dmy0  xr0_4__dmy0 xr0_5__dmy0  rppolyhri3d3k lr=7.34e-6 wr=2e-6 mf=1 m=1 mismatchflag=1
xr0_6__dmy0  xr0_5__dmy0 net029  rppolyhri3d3k lr=7.34e-6 wr=2e-6 mf=1 m=1 mismatchflag=1

.ENDS
