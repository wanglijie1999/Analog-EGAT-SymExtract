** Generated for: hspiceD
** Generated on: Mar  9 09:51:24 2023
** Design library name: DDA_22Train
** Design cell name: DDA_2021_MQQ
** Design view name: schematic



** Library name: DDA_22Train
** Cell name: DDA_2021_MQQ
** View name: schematic
.subckt 05DDAMQQ vss vo vdd ibias _net0 _net1 _net2 _net3
xm29 vss vss vss vss nch_5 l=2e-6 w=2e-6 m=30 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm6 net45 vb net39 vss nch_5 l=2e-6 w=2e-6 m=6 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm0 ibias ibias net47 vss nch_5 l=2e-6 w=2e-6 m=1 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm5 net29 net29 vss vss nch_5 l=2e-6 w=2e-6 m=4 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm4 net65 net47 vss vss nch_5 l=2e-6 w=2e-6 m=2 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm3 net47 net47 vss vss nch_5 l=2e-6 w=2e-6 m=1 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm2 vb vb net29 vss nch_5 l=2e-6 w=2e-6 m=4 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm7 vo vb net36 vss nch_5 l=2e-6 w=2e-6 m=6 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm1 net33 ibias net65 vss nch_5 l=2e-6 w=2e-6 m=2 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm8 net39 net47 vss vss nch_5 l=2e-6 w=2e-6 m=10 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm9 net36 net47 vss vss nch_5 l=2e-6 w=2e-6 m=10 nf=1 sd=540e-9 ad=960e-15 as=960e-15 pd=4.96e-6 ps=4.96e-6 nrd=135e-3 nrs=135e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm28 vdd vdd vdd vdd pch_5 l=1e-6 w=4e-6 m=8 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm27 net033 net033 net033 net033 pch_5 l=1e-6 w=8e-6 m=4 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm26 net025 net025 net025 net025 pch_5 l=1e-6 w=8e-6 m=4 nf=1 sd=540e-9 ad=3.84e-12 as=3.84e-12 pd=16.96e-6 ps=16.96e-6 nrd=33.75e-3 nrs=33.75e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm22 net45 net45 net46 vdd pch_5 l=1e-6 w=4e-6 m=6 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm21 net39 _net2 net033 net033 pch_5 l=2e-6 w=32e-6 m=2 nf=4 sd=540e-9 ad=8.64e-12 as=12e-12 pd=34.16e-6 ps=51e-6 nrd=8.4375e-3 nrs=8.4375e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm16 net36 _net0 net025 net025 pch_5 l=2e-6 w=32e-6 m=2 nf=4 sd=540e-9 ad=8.64e-12 as=12e-12 pd=34.16e-6 ps=51e-6 nrd=8.4375e-3 nrs=8.4375e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm12 net64 net34 vdd vdd pch_5 l=1e-6 w=4e-6 m=1 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm17 net39 _net1 net025 net025 pch_5 l=2e-6 w=32e-6 m=2 nf=4 sd=540e-9 ad=8.64e-12 as=12e-12 pd=34.16e-6 ps=51e-6 nrd=8.4375e-3 nrs=8.4375e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm18 net61 net34 vdd vdd pch_5 l=1e-6 w=4e-6 m=5 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm24 vo net45 net63 vdd pch_5 l=1e-6 w=4e-6 m=6 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm15 net025 net33 net62 vdd pch_5 l=1e-6 w=4e-6 m=5 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm11 vb net33 net64 vdd pch_5 l=1e-6 w=4e-6 m=1 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm20 net36 _net3 net033 net033 pch_5 l=2e-6 w=32e-6 m=2 nf=4 sd=540e-9 ad=8.64e-12 as=12e-12 pd=34.16e-6 ps=51e-6 nrd=8.4375e-3 nrs=8.4375e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm19 net033 net33 net61 vdd pch_5 l=1e-6 w=4e-6 m=5 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm14 net62 net34 vdd vdd pch_5 l=1e-6 w=4e-6 m=5 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm10 net33 net33 net34 vdd pch_5 l=1e-6 w=4e-6 m=2 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm23 net46 net46 vdd vdd pch_5 l=1e-6 w=4e-6 m=4 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm25 net63 net46 vdd vdd pch_5 l=1e-6 w=4e-6 m=4 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
xm13 net34 net34 vdd vdd pch_5 l=1e-6 w=4e-6 m=2 nf=1 sd=540e-9 ad=1.92e-12 as=1.92e-12 pd=8.96e-6 ps=8.96e-6 nrd=67.5e-3 nrs=67.5e-3 sa=480e-9 sb=480e-9 sca=0 scb=0 scc=0
.ENDS
